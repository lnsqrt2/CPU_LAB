#include "stdi.v"
module test()
wire;
reg test[1:0];

endmodule