
module divider(clk_in, clk_out)

input clk_in;
output clk_out;

reg clk_out;

endmodule