module regfile()
wire;
reg test[1:0];

endmodule